LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
ENTITY MUX21A2130 IS
	
	PORT(a,b:IN STD_LOGIC;
			 s:IN STD_LOGIC;
          y:OUT STD_LOGIC);
			 
END ENTITY MUX21A2130;

ARCHITECTURE one OF MUX21A2130 IS BEGIN 
	PROCESS (a,b,s) BEGIN
		IF S = '0' THEN
			y <= a;
		ELSE
			y <= b;
		END IF;
	END PROCESS;
END ARCHITECTURE ONE;